module app

@[heap]
pub struct Session {
	pub mut:
	is_open       bool
}
