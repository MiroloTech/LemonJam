module uilib

@[heap]
pub struct ParticleEmitter {
	pub mut:
	amount              int            = 20
	seperate_draw_call  bool           = true
	// TODO : This ( just for fun and more app juice )
}
