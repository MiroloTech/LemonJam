module objs

pub struct Instrument {
	pub mut:
	name         string
	icon         string
}
