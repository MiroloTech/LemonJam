module objs

pub struct Effect {
	pub mut:
	name         string
	icon         string
}
