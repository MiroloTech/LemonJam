module mirrorlib

// List of basic action codes for easier use

pub const action_user_connected                := u32(0)
pub const action_join_session_hash             := u32(1)
pub const action_heartbeat                     := u32(2)
pub const action_lock_nid                      := u32(3)
pub const action_unlock_nid                    := u32(4)
