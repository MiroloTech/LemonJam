module objs

pub struct Pattern {
	pub mut:
	name         string
	notes        []&Note
}

